// module tb2;

// reg [6:0] address;
// wire [31:0] instruction;

// instructionMemory im(instruction, address);


// initial
// 	begin
// // 		$monitor("%t %b %b", $time, address, instruction);
// // 		# 5 address <= 6'b000000;
// // 		# 10 address <= 6'b000001;
// // 		# 15 address <= 6'b000010;
// // 		# 20 address <= 6'b000011;
		
// // 		# 100000 $finish;
// 	end

// endmodule
