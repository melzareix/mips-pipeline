// module tb5;
// reg [31:0] reg1,reg2;
// reg [2:0] ALUcontrol;
 
// wire [31:0] out;
// wire zeroFlag;
// ALU A(zeroFlag,out,reg1,reg2,ALUcontrol);
 


//  initial
//  begin  
//  fork
//  		// $monitor("%t %b %b", $time, out,zeroFlag);
//    //      # 5 reg1 <= 32'b00000111011111111101111111111111; reg2 <= 32'b00000111011111111101111111111111; 
//    //      # 10 ALUcontrol <= 3'b000;
//    //      # 15 ALUcontrol <= 3'b001;
//    //      # 20 ALUcontrol <= 3'b010;
//    //      # 25 ALUcontrol <= 3'b011;
//    //      # 30 ALUcontrol <= 3'b100;
//    //      # 35 ALUcontrol <= 3'b101;
//    //      # 40 ALUcontrol <= 3'b011;
//    //      # 45 reg2<= 32'b11111111111111111111111111111111;
//    //      # 50 ALUcontrol <= 3'b101;
//    //      # 55 ALUcontrol <= 3'b110;
//    //      # 60 reg1 <= 32'b1;
//    //      # 65 reg2<= 32'b0;
        
        
//    //  	# 65 $finish;
// join
//  end
 

// endmodule
