
module Processor_tb;


Processor r();
endmodule